`ifndef CONST_VH
`define CONST_VH
`define HTIF_WIDTH 16
`define MEM_DATA_BITS 128
`define buffer_sram false
`define MEM_TAG_BITS 6
`define MEM_ADDR_BITS 26
`endif // CONST_VH
